import rv32i_types::*;

module load_store_q
(
	input sal_t rob_bus,
	input rs_t rs1_out,
	input 
);


endmodule : load_store_q
