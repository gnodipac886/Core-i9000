module l2_cache_control #(parameter NUM_WAYS = 8,
                        parameter WAYS_LOG_2 = $clog2(NUM_WAYS))
(
  input clk,

  /* CPU memory data signals */
  input  logic mem_read,
	input  logic mem_write,
	output logic mem_resp,

  /* Physical memory data signals */
  input  logic pmem_resp,
	output logic pmem_read,
	output logic pmem_write,

  /* Control signals */
  output logic tag_load,
  output logic valid_load,
  output logic dirty_load,
  output logic dirty_in,
  input logic dirty_out,

  input logic hit,
  output logic [1:0] writing,

  input logic [WAYS_LOG_2 - 1:0] lru_out[NUM_WAYS],
  input logic [WAYS_LOG_2 - 1 : 0] _idx,
  input logic valid_out[NUM_WAYS],
  output logic lru_load[NUM_WAYS],
  output logic [WAYS_LOG_2 - 1:0] lru_in [NUM_WAYS]
);

/* State Enumeration */
enum int unsigned
{
  check_hit,
	read_mem
} state, next_state;

//          0 1 2 3 4 5 6 7
// valid:   1 0 0 0 0 0 0 0
// lru:     0 7 7 7 7 7 7 7

function void update_lru();
  for (int i = 0; i < NUM_WAYS; i++ ) begin
    if (valid_out[i] && (lru_out[i] < lru_out[_idx])) begin
      lru_load[i] = 1'b1;
      lru_in[i] = lru_out[i] + 1;
    end
  end
  lru_load[_idx] = 1'b1;
  lru_in[_idx] = '0;
endfunction

/* State Control Signals */
always_comb begin : state_actions

	/* Defaults */
  tag_load = 1'b0;
  valid_load = 1'b0;
  dirty_load = 1'b0;
  dirty_in = 1'b0;
  writing = 2'b11;

	mem_resp = 1'b0;
	pmem_write = 1'b0;
	pmem_read = 1'b0;

  for(int i = 0; i < NUM_WAYS; i++) begin 
    lru_load[i] = 1'b0;
    lru_in[i] = 0;
  end 

	case(state)
    check_hit: begin
      if (mem_read || mem_write) begin
        if (hit) begin
          mem_resp = 1'b1;
          if (mem_write) begin
            dirty_load = 1'b1;
            dirty_in = 1'b1;
            writing = 2'b01;
          end
          update_lru();
        end else begin
          if (dirty_out)
            pmem_write = 1'b1;
        end
      end
    end

    read_mem: begin
      pmem_read = 1'b1;
      writing = 2'b00;
      if (pmem_resp) begin
        tag_load = 1'b1;
        valid_load = 1'b1;
      end
        dirty_load = 1'b1;
        dirty_in = 1'b0;
    end

	endcase
end

/* Next State Logic */
always_comb begin : next_state_logic

	/* Default state transition */
	next_state = state;

	case(state)
    check_hit: begin
      if ((mem_read || mem_write) && !hit) begin
        if (dirty_out) begin
          if (pmem_resp)
            next_state = read_mem;
        end else begin
          next_state = read_mem;
		  end
      end
    end

    read_mem: begin
      if (pmem_resp)
        next_state = check_hit;
    end

	endcase
end

/* Next State Assignment */
always_ff @(posedge clk) begin: next_state_assignment
	 state <= next_state;
end

endmodule : l2_cache_control
