import rv32i_types::*;

module load_store_q
(
	
);


endmodule : load_store_q
