module fetcher #(parameter width = 32)
(
	input clk,
	input rst,
	input dequeue,
	input [width-1:0] in,
	output logic [width-1:0] out
);


	register MDR(
		.load(),
		.in(),
		.out(),
		.*
	);

endmodule : fetcher
